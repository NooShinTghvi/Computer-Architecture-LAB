module IF (
		input clk,rst,freez, BrTaken,
		// SRAM  UNIT
		pause,
		input [31:0] BrAdder, output [31:0] PC,instruction
	);

	wire [31:0] PCIn,instructionIn;

	IFSub _IFsub (clk,rst,freez,BrTaken,pause,BrAdder,PCIn,instructionIn);
	IFReg _IFReg (clk,rst,freez, BrTaken,pause, PCIn,instructionIn,PC,instruction);

endmodule

// * * * * * * * * * * * * * * * * * * * * * * * * * * * * * * * *
module IFSub (input clk,rst,freez,BrTaken,pause,input [31:0] BrAdder, output [31:0] PC4,output [31:0] Instruction);
	reg [31:0] ram [1023:0]; //2 ^ 10 = 1024
	wire [31:0] PCMuxOut;
	reg [31:0] PC; //
	integer i;
	initial begin
		ram[0] = 32'b10000000000000010000011000001010;//-- Addi r1 ,r0 ,1546
		ram[4] = 32'b00000100000000010001000000000000;//-- Add  r2 ,r0 ,r1
		ram[8] = 32'b00001100000000010001100000000000;//-- sub r3 ,r0 ,r1
		ram[12] = 32'b00010100010000110010000000000000;//-- And r4 ,r2 ,r3
		ram[16] = 32'b10000100011001010001101000110100;//-- Subi r5 ,r3 ,6708
		ram[20] = 32'b00011000011001000010100000000000;//-- or r5 ,r3 ,r4
		ram[24] = 32'b00011100101000000011000000000000;//-- nor  r6 ,r5 ,r0
		ram[28] = 32'b00011100100000000101100000000000;//-- nor  r11 ,r4 ,r0
		ram[32] = 32'b00001100101001010010100000000000;//-- sub r5 ,r5 ,r5
		ram[36] = 32'b10000000000000010000010000000000;//-- Addi  r1 ,r0 ,1024 ** 10
		ram[40] = 32'b10010100001000100000000000000000;//-- st r2 ,r1 ,0
		ram[44] = 32'b10010000001001010000000000000000;//-- ld r5 ,r1 ,0
		ram[48] = 32'b10100000101000000000000000000001;//-- Bez r5 ,1
		ram[52] = 32'b00100000101000010011100000000000;//-- xor r7 ,r5 ,r1
		ram[56] = 32'b00100000101000010000000000000000;//-- xor r0 ,r5 ,r1
		ram[60] = 32'b00100100011010110011100000000000;//-- sla r7 ,r3 ,r11
		ram[64] = 32'b00101000011010110100000000000000;//-- sll r8 ,r3 ,r11
		ram[68] = 32'b00101100011001000100100000000000;//-- sra r9 ,r3 ,r4
		ram[72] = 32'b00110000011001000101000000000000;//-- srl r10 ,r3 ,r4
		ram[76] = 32'b10010100001000110000000000000100;//-- st r3 ,r1 ,4  **20
		ram[80] = 32'b10010100001001000000000000001000;//-- st r4 ,r1 ,8
		ram[84] = 32'b10010100001001010000000000001100;//-- st r5 ,r1 ,12
		ram[88] = 32'b10010100001001100000000000010000;//-- st r6 ,r1 ,16
		ram[92] = 32'b10010000001010110000000000000100;//-- ld r11 ,r1 ,4 wite? miss
		ram[96] = 32'b10010100001001110000000000010100;//-- st r7 ,r1 ,20
		ram[100] = 32'b10010100001010000000000000011000;//-- st r8 ,r1 ,24
		ram[104] = 32'b10010100001010010000000000011100;//-- st r9 ,r1 ,28
		ram[108] = 32'b10010100001010100000000000100000;//-- st r10 ,r1 ,32
		ram[112] = 32'b10010100001010110000000000100100;//-- st r11 ,r1 ,36
		ram[116] = 32'b10000000000000010000000000000011;//-- Addi  r1 ,r0 ,3 **30
		ram[120] = 32'b10000000000001000000010000000000;//-- Addi r4 ,r0 ,1024
		ram[124] = 32'b10000000000000100000000000000000;//-- Addi  r2 ,r0 ,0
		ram[128] = 32'b10000000000000110000000000000001;//-- Addi  r3 ,x ,1   <--- Jump 2
		ram[132] = 32'b10000000000010010000000000000010;//-- Addi  r9 ,r0 ,2   <--- Jump 1
		ram[136] = 32'b00101000011010010100000000000000;//-- sll r8 ,r3 ,r9
		ram[140] = 32'b00000100100010000100000000000000;//-- Add  r8 ,r4 ,r8
		ram[144] = 32'b10010001000001010000000000000000;//-- ld r5 ,r8 ,0 //hit
		ram[148] = 32'b10010001000001101111111111111100;//-- ld r6 ,r8 ,-4
		ram[152] = 32'b00001100101001100100100000000000;//-- sub  r9 ,r5 ,r6
		ram[156] = 32'b10000000000010101000000000000000;//-- Addi  r10 ,r0 ,0x8000 **40
		ram[160] = 32'b10000000000010110000000000010000;//-- Addi r11 ,r0 ,16
		ram[164] = 32'b00101001010010110101000000000000;//-- sll r10 ,r1 ,r11
		ram[168] = 32'b00010101001010100100100000000000;//-- And  r9 ,r9 ,r10
		ram[172] = 32'b10100001001000000000000000001000;//-- Bez r9 ,4
		ram[176] = 32'b100101_01000_00101_1111111111111100;//-- st r5 ,r8 ,-4
		ram[180] = 32'b100101_01000_00110_0000000000000000;//-- st r6 ,r8 ,0
		ram[184] = 32'b100000_00011_00011_0000000000000001;//-- Addi  r3 ,r3 ,1
		ram[188] = 32'b101001_00001_00011_1111111111000100;//-- BNE r1 ,r3 ,-15 ---> Jump 1
		ram[192] = 32'b10000000010000100000000000000001;//-- Addi  r2 ,r2 ,1
		ram[196] = 32'b10100100001000101111111110111000;//-- BNE r1 ,r2 ,-18 **50  ----> Jump 2
		ram[200] = 32'b10000000000000010000010000000000;//-- Addi  r1 ,r0 ,1024
		ram[204] = 32'b10010000001000100000000000000000;//-- ld ,r2 ,r1 ,0
		ram[208] = 32'b10010000001000110000000000000100;//-- ld ,r3 ,r1 ,4
		ram[212] = 32'b10010000001001000000000000001000;//-- ld ,r4 ,r1 ,8
		ram[216] = 32'b10010000001001000000001000001000;//-- ld ,r4 ,r1 ,520
		ram[220] = 32'b10010000001001000000010000001000;//-- ld ,r4 ,r1 ,1023
		ram[224] = 32'b10010000001001010000000000001100;//-- ld ,r5 ,r1 ,12
		ram[228] = 32'b10010000001001100000000000010000;//-- ld ,r6 ,r1 ,16
		ram[232] = 32'b10010000001001110000000000010100;//-- ld ,r7 ,r1 ,20
		ram[236] = 32'b10010000001010000000000000011000;//-- ld ,r8 ,r1 ,24 **60
		ram[240] = 32'b10010000001010010000000000011100;//-- ld ,r9 ,r1 ,28
		ram[244] = 32'b10010000001010100000000000100000;//-- ld ,r10,r1 ,32
		ram[248] = 32'b10010000001010110000000000100100;//-- ld ,r11,r1 ,36
		ram[252] = 32'b10101000000000001111111111111100;//-- JMP  -1 **64
	end

	assign PC4 = PC + 4;	// PC + 4

	Mux2to1_32 _PCBrMux(BrTaken,PC4,BrAdder,PCMuxOut);

	always@(posedge clk,posedge rst) begin //Read from ram
		if (rst) begin
			PC = 32'd0;
		end
		else begin
			if (freez == 1'b1 || pause == 1'b1) begin
				PC = PC;
			end
			else begin
				PC = PCMuxOut;
			end
		end
	end
	assign Instruction = ram[{PC[31:2],2'b0}];

endmodule
// * * * * * * * * * * * * * * * * * * * * * * * * * * * * * * * *

module IFReg (
		input clk,rst,freez, BrTaken,
		// SRAM  UNIT
		pause,
		input[31:0] PCin,instructionIn,output reg [31:0] PC,instruction
	);
	always@(posedge clk,posedge rst) begin
		if (rst) begin
			PC <= 32'd0;
			instruction <= 32'd0;
		end
		else if(BrTaken)
			instruction <= 32'b0;
		else begin
			if (freez == 1'b1 || pause == 1'b1) begin
				PC <= PC;
				instruction <= instruction;
			end
			else begin
				PC <= PCin;
				instruction <= instructionIn;
			end
		end
	end
endmodule
// * * * * * * * * * * * * * * * * * * * * * * * * * * * * * * * *
